module mul(input [7:0] mc, input [7:0] mp, output [15:0] p);
    assign p = mc * mp;
endmodule
